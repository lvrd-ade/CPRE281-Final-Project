module mux8to1 (
    input [7:0] w0, w1, w2, w3, w4, w5, w6, w7,
    input [2:0] s,
    output reg [7:0] f
);
always @(*)
begin
    case(s)
        3'b000: f = w0;
        3'b001: f = w1;
        3'b010: f = w2;
        3'b011: f = w3;
        3'b100: f = w4;
        3'b101: f = w5;
        3'b110: f = w6;
        3'b111: f = w7;
    endcase
end
endmodule
